../bsg_repo/bsg_misc/bsg_counter_clear_up.sv