../bsg_repo/bsg_misc/bsg_defines.sv