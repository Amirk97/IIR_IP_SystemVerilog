module IIR

  endmodule
